module sig_cntrl (opcode,opcode_ext,reg2_rd_sel, jump, im_sel, ALU_src, wb_sel, wb_sel0, wb_sel1, ex_result_sel, invRs, invIn, Cin, ALUOP, alu_sign, MemWrite, MemRead, reg_write,Branch_op, rd_sel, mem_en, BranchEn,
		JumpReg, Halt, s_extend, LBI_sel, SLBI_sel, BTR_sel, STU_sel, isBranch, Read1, Read2, write_from_mem, wreg_flag, isJR);
    input [4:0] opcode;
	input [1:0] opcode_ext;
    output reg reg2_rd_sel, jump, im_sel, ALU_src, wb_sel, wb_sel1, ex_result_sel, invRs, invIn, Cin, alu_sign, MemWrite, MemRead, reg_write, mem_en, BranchEn, JumpReg, s_extend, LBI_sel, SLBI_sel, BTR_sel, STU_sel,
				isBranch, Read1, Read2, write_from_mem, wreg_flag, isJR;
    output Halt;
	output reg [1:0] Branch_op, rd_sel, wb_sel0;
	output reg [2:0] ALUOP;

	assign Halt = & (~ opcode[4:0]);

always @ (*) begin
    case(opcode)
		5'b00001:  begin    //NOP
			reg_write <= 1'b0;
			reg2_rd_sel <= 1'b0;
			im_sel <= 1'b0;
			rd_sel <= 2'b01;
			ALU_src <= 1'b0;
			jump <= 1'b0;
			MemWrite <= 1'b0;
			MemRead <= 1'b0;
			wb_sel <= 1'b1;
			wb_sel0 <= 2'b00;
			wb_sel1 <= 1'b0;
			ex_result_sel <= 1'b1;
			s_extend <= 1;
			invRs <= 1'b0;
			invIn <= 1'b0;
			Cin <= 1'b0;
			ALUOP <= 3'b100;
			alu_sign<= 1'b1;
			Branch_op <= 2'b00;
			mem_en <= 1'b0;
			BranchEn <= 1'b0;
			JumpReg <= 1'b0;
			LBI_sel <= 1'b0;
			SLBI_sel <= 1'b0;
			BTR_sel <= 1'b0;
			STU_sel <= 1'b0;
			isBranch <= 1'b0;
			Read1 <= 1'b0;
			Read2 <= 1'b0;
			write_from_mem <= 1'b0;
			wreg_flag <= 1'b0;
			isJR <= 1'b0;
		end
	    5'b01000:  begin    //ADDI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b100;
				alu_sign<= 1'b1;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b01001:  begin // SUBI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b1;
				invIn <= 1'b0;
				Cin <= 1'b1;
				ALUOP <= 3'b100;
				alu_sign<= 1'b1;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b01010:  begin  // XORI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 0;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b111;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b01011:  begin // ANDNI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 0;
				invRs <= 1'b0;
				invIn <= 1'b1;
				Cin <= 1'b0;
				ALUOP <= 3'b101;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10100:  begin  // ROLI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b000;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10101:  begin  // SLLI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b001;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10110:  begin  // RORI Rd, Rs, immediate R
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b010;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10111:  begin  // SRLI Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b011;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10000:  begin  // ST Rd, Rs, immediate
		        reg_write <= 1'b0;
				reg2_rd_sel <= 1'b1;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b1;
				MemRead <= 1'b0;
				wb_sel <= 1'b0;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b100;
				alu_sign<= 1'b1;
				Branch_op <= 2'b00;
				mem_en <= 1'b1;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b1;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
            end
		5'b10001:  begin  // LD Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b1;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b1;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b100;
				alu_sign<= 1'b1;
				Branch_op <= 2'b00;
				mem_en <= 1'b1;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b1;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10011:  begin  // STU Rd, Rs, immediate
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b1;
				im_sel <= 1'b0;
				rd_sel <= 2'b01;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b1;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 3'b100;
				alu_sign<= 1'b1;
				Branch_op <= 2'b00;
				mem_en <= 1'b1;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b0;
				STU_sel <= 1'b1;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b1;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b11001:  begin  // BTR Rd, Rs
		        reg_write <= 1'b1;
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b00;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0;
				MemRead <= 1'b0;
				wb_sel <= 1'b1;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				s_extend <= 1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 1'b0;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 1'b0;
				SLBI_sel <= 1'b0;
				BTR_sel <= 1'b1;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b11011:  begin
				case (opcode_ext)
				2'b00: begin  // ADD Rd, Rs, Rt
					reg_write <= 1'b1;
					reg2_rd_sel <= 1'b0;
					im_sel <= 1'b0;
					rd_sel <= 2'b00;
					ALU_src <= 1'b1;
					jump <= 1'b0;
					MemWrite <= 1'b0;
					MemRead <= 1'b0;
					wb_sel <= 1'b1;
					wb_sel0 <= 2'b00;
					wb_sel1 <= 1'b0;
					ex_result_sel <= 1'b1;
					s_extend <= 1;
					invRs <= 1'b0;
					invIn <= 1'b0;
					Cin <= 1'b0;
					ALUOP <= 3'b100;
					alu_sign<= 1'b0;
					Branch_op <= 2'b00;
					mem_en <= 1'b0;
					BranchEn <= 1'b0;
					JumpReg <= 1'b0;
					LBI_sel <= 1'b0;
					SLBI_sel <= 1'b0;
					BTR_sel <= 1'b0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
						end
				2'b01: begin // SUB Rd, Rs, Rt
					reg_write <= 1'b1;
					reg2_rd_sel <= 1'b0;
					im_sel <= 1'b0;
					rd_sel <= 2'b00;
					ALU_src <= 1'b1;
					jump <= 1'b0;
					MemWrite <= 1'b0;
					MemRead <= 1'b0;
					wb_sel <= 1'b1;
					wb_sel0 <= 2'b00;
					wb_sel1 <= 1'b0;
					ex_result_sel <= 1'b1;
					s_extend <= 1;
					invRs <= 1'b1;
					invIn <= 1'b0;
					Cin <= 1'b1; // 2's complement must add 1
					ALUOP <= 3'b100;
					alu_sign<= 1'b0;
					Branch_op <= 2'b00;
					mem_en <= 1'b0;
					BranchEn <= 1'b0;
					JumpReg <= 1'b0;
					LBI_sel <= 1'b0;
					SLBI_sel <= 1'b0;
					BTR_sel <= 1'b0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
				        end
				2'b10: begin // XOR Rd, Rs, Rt
					reg_write <= 1'b1;
					reg2_rd_sel <= 1'b0;
					im_sel <= 1'b0;
					rd_sel <= 2'b00;
					ALU_src <= 1'b1;
					jump <= 1'b0;
					MemWrite <= 1'b0;
					MemRead <= 1'b0;
					wb_sel <= 1'b1;
					wb_sel0 <= 2'b00;
					wb_sel1 <= 1'b0;
					ex_result_sel <= 1'b1;
					s_extend <= 1;
					invRs <= 1'b0;
					invIn <= 1'b0;
					Cin <= 1'b0;
					ALUOP <= 3'b111;
					alu_sign<= 1'b0;
					Branch_op <= 2'b00;
					mem_en <= 1'b0;
					BranchEn <= 1'b0;
					JumpReg <= 1'b0;
					LBI_sel <= 1'b0;
					SLBI_sel <= 1'b0;
					BTR_sel <= 1'b0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
						end
				2'b11: begin // ANDN Rd, Rs, Rt
					reg_write <= 1'b1;
					reg2_rd_sel <= 1'b0;
					im_sel <= 1'b0;
					rd_sel <= 2'b00;
					ALU_src <= 1'b1;
					jump <= 1'b0;
					MemWrite <= 1'b0;
					MemRead <= 1'b0;
					wb_sel <= 1'b1;
					wb_sel0 <= 2'b00;
					wb_sel1 <= 1'b0;
					ex_result_sel <= 1'b1;
					s_extend <= 1;
					invRs <= 1'b0;
					invIn <= 1'b1;
					Cin <= 1'b0;
					ALUOP <= 3'b101;
					alu_sign<= 1'b0;
					Branch_op <= 2'b00;
					mem_en <= 1'b0;
					BranchEn <= 1'b0;
					JumpReg <= 1'b0;
					LBI_sel <= 1'b0;
					SLBI_sel <= 1'b0;
					BTR_sel <= 1'b0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
				end
				endcase
            end

	5'b11010:  begin
			case (opcode_ext)
				2'b00: begin  // ROL Rd, Rs, Rt
					reg2_rd_sel <= 0;
					jump <= 0;
					im_sel <= 0;
					ALU_src <= 1;
					wb_sel <= 1;
					wb_sel0 <= 0;
					wb_sel1 <= 0;
					ex_result_sel <= 1'b1;
					invRs <= 0;
					invIn <= 0;
					Cin <= 0;
					ALUOP <= 0;
					alu_sign <= 0;
					MemWrite <= 0;
					MemRead <= 1'b0;
					reg_write <= 1;
					Branch_op <= 0;
					rd_sel <= 0;
					mem_en <= 0;
					BranchEn <= 0;
					JumpReg <= 0;
					s_extend <= 1;
					LBI_sel <= 0;
					SLBI_sel <= 0;
					BTR_sel <= 0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
					end
				2'b01: begin // SLL Rd, Rs, Rt
					reg2_rd_sel <= 0;
					jump <= 0;
					im_sel <= 0;
					ALU_src <= 1;
					wb_sel <= 1;
					wb_sel0 <= 0;
					wb_sel1 <= 0;
					ex_result_sel <= 1'b1;
					invRs <= 0;
					invIn <= 0;
					Cin <= 0;
					ALUOP <= 1;
					alu_sign <= 0;
					MemWrite <= 0;
					MemRead <= 1'b0;
					reg_write <= 1;
					Branch_op <= 0;
					rd_sel <= 0;
					mem_en <= 0;
					BranchEn <= 0;
					JumpReg <= 0;
					s_extend <= 1;
					LBI_sel <= 0;
					SLBI_sel <= 0;
					BTR_sel <= 0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
					end
				2'b10: begin  // ROR Rd, Rs, Rt
					reg2_rd_sel <= 0;
					jump <= 0;
					im_sel <= 0;
					ALU_src <= 1;
					wb_sel <= 1;
					wb_sel0 <= 0;
					wb_sel1 <= 0;
					ex_result_sel <= 1'b1;
					invRs <= 0;
					invIn <= 0;
					Cin <= 0;
					ALUOP <= 2;
					alu_sign <= 0;
					MemWrite <= 0;
					MemRead <= 1'b0;
					reg_write <= 1;
					Branch_op <= 0;
					rd_sel <= 0;
					mem_en <= 0;
					BranchEn <= 0;
					JumpReg <= 0;
					s_extend <= 1;
					LBI_sel <= 0;
					SLBI_sel <= 0;
					BTR_sel <= 0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
					end
				2'b11: begin //SRL Rd, Rs, Rt
					reg2_rd_sel <= 0;
					jump <= 0;
					im_sel <= 0;
					ALU_src <= 1;
					wb_sel <= 1;
					wb_sel0 <= 0;
					wb_sel1 <= 0;
					ex_result_sel <= 1'b1;
					invRs <= 0;
					invIn <= 0;
					Cin <= 0;
					ALUOP <= 3;
					alu_sign <= 0;
					MemWrite <= 0;
					MemRead <= 1'b0;
					reg_write <= 1;
					Branch_op <= 0;
					rd_sel <= 0;
					mem_en <= 0;
					BranchEn <= 0;
					JumpReg <= 0;
					s_extend <= 1;
					LBI_sel <= 0;
					SLBI_sel <= 0;
					BTR_sel <= 0;
					STU_sel <= 1'b0;
					isBranch <= 1'b0;
					Read1 <= 1'b1;
					Read2 <= 1'b1;
					write_from_mem <= 1'b0;
					wreg_flag <= 1'b1;
					isJR <= 1'b0;
					end
				default: begin
					reg2_rd_sel <= 0;
					jump <= 0;
					im_sel <= 0;
					ALU_src <= 0;
					wb_sel <= 0;
					wb_sel0 <= 0;
					wb_sel1 <= 0;
					ex_result_sel <= 1'b1;
					invRs <= 0;
					invIn <= 0;
					Cin <= 0;
					ALUOP <= 0;
					alu_sign <= 0;
					MemWrite <= 0;
					MemRead <= 1'b0;
					reg_write <= 0;
					Branch_op <= 0;
					rd_sel <= 0;
					mem_en <= 0;
					BranchEn <= 0;
					JumpReg <= 0;
					s_extend <= 1;
					LBI_sel <= 0;
					SLBI_sel <= 0;
					BTR_sel <= 0;
					STU_sel <= 1'b0;
					isJR <= 1'b0;
					end
				endcase
            end
		5'b11100:  begin  // SEQ Rd, Rs, Rt
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 0;
				ALU_src <= 1;
				wb_sel <= 1;
				wb_sel0 <= 2;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b0;
				invRs <= 0;
				invIn <= 1;
				Cin <= 1;
				ALUOP <= 4;
				alu_sign <= 1;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b1;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b11101:  begin  // SLT Rd, Rs, Rt
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 0;
				ALU_src <= 1;
				wb_sel <= 1;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b0;
				invRs <= 0;
				invIn <= 1;
				Cin <= 1;
				ALUOP <= 4;
				alu_sign <= 1;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b1;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b11110:  begin  // SLE Rd, Rs, Rt
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 0;
				ALU_src <= 1;
				wb_sel <= 1;
				wb_sel0 <= 1;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b0;
				invRs <= 0;
				invIn <= 1;
				Cin <= 1;
				ALUOP <= 4;
				alu_sign <= 1;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b1;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b11111:  begin  //SCO Rd, Rs, Rt
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 0;
				ALU_src <= 1;
				wb_sel <= 1;
				wb_sel0 <= 3;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b0;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 4;
				alu_sign <= 1;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b1;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b01100:  begin  // BEQZ Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 0;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 1;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b1;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
            end
		5'b01101:  begin  //BNEZ Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 0;
				Branch_op <= 1;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 1;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b1;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
            end
		5'b01110:  begin  //BLTZ Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 0;
				Branch_op <= 2;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 1;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b1;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
            end
		5'b01111:  begin  //BGEZ Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 0;
				Branch_op <= 3;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 1;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b1;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
            end
		5'b11000:  begin  // LBI Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 2;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 1;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b0;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b10010:  begin  //SLBI Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 1;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 6;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 2;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 0;
				LBI_sel <= 0;
				SLBI_sel <= 1;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b00100:  begin  //J displacement
				reg2_rd_sel <= 0;
				jump <= 1;
				im_sel <= 0;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 0;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b1;
				Read1 <= 1'b0;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
            end
		5'b00101:  begin   //JR Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 4;
				alu_sign <= 1;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 0;
				Branch_op <= 0;
				rd_sel <= 0;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 1;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b1;
            end
		5'b00110:  begin  //JAL displacement
				reg2_rd_sel <= 0;
				jump <= 1;
				im_sel <= 0;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 0;
				alu_sign <= 0;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 3;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 0;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b1;
				Read1 <= 1'b0;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b0;
            end
		5'b00111:  begin  //JALR Rs, immediate
				reg2_rd_sel <= 0;
				jump <= 0;
				im_sel <= 1;
				ALU_src <= 0;
				wb_sel <= 0;
				wb_sel0 <= 0;
				wb_sel1 <= 0;
				ex_result_sel <= 1'b1;
				invRs <= 0;
				invIn <= 0;
				Cin <= 0;
				ALUOP <= 4;
				alu_sign <= 1;
				MemWrite <= 0;
				MemRead <= 1'b0;
				reg_write <= 1;
				Branch_op <= 0;
				rd_sel <= 3;
				mem_en <= 0;
				BranchEn <= 0;
				JumpReg <= 1;
				s_extend <= 1;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b1;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b1;
				isJR <= 1'b1;
            end
		default: begin
				reg_write <= 1'b0; //always 0 at default
				reg2_rd_sel <= 1'b0;
				im_sel <= 1'b0;
				rd_sel <= 2'b00;
				ALU_src <= 1'b0;
				jump <= 1'b0;
				MemWrite <= 1'b0; //always 0 at default
				MemRead <= 1'b0;
				wb_sel <= 1'b0;
				wb_sel0 <= 2'b00;
				wb_sel1 <= 1'b0;
				ex_result_sel <= 1'b1;
				invRs <= 1'b0;
				invIn <= 1'b0;
				Cin <= 1'b0;
				ALUOP <= 1'b0;
				alu_sign<= 1'b0;
				Branch_op <= 2'b00;
				rd_sel <= 2'b00;
				mem_en <= 1'b0;
				BranchEn <= 1'b0;
				JumpReg <= 1'b0;
				LBI_sel <= 0;
				SLBI_sel <= 0;
				BTR_sel <= 0;
				STU_sel <= 1'b0;
				isBranch <= 1'b0;
				Read1 <= 1'b0;
				Read2 <= 1'b0;
				write_from_mem <= 1'b0;
				wreg_flag <= 1'b0;
				isJR <= 1'b0;
				end
	endcase
end
endmodule
